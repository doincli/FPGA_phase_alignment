    .INIT_00(256'h0000000ba252f03200000001b000100100000020a4f2f01e00000020a3101000),
    .INIT_01(256'h00000014a00206dc0000000ba26206e000000014b002070000000014a0e20767),
    .INIT_02(256'h00000014a002b20f00000014b002089400000014a00206da00000014b0022478),
    .INIT_03(256'h0000002f21d2f032000000062b0010020000000b21d2b80f00000014b002b40f),
    .INIT_04(256'h00000014b00206dc00000014a002071400000014b00224b900000014a0020767),
    .INIT_05(256'h00000014b00206b400000014a000bc0a00000014b00206b400000014a000bc0b),
    .INIT_06(256'h00000014a00206b40000000ba270bc0800000014b00206b400000014a000bc09),
    .INIT_07(256'h00000014a000900200000014b00206da00000014a00206b400000014b000bc07),
    .INIT_08(256'h0000002fb1c0101000000006b20208940000000b21c3242600000014b000d008),
    .INIT_09(256'h0000000d1ff2074b00000001b000100000000001a0022008000000250002074b),
    .INIT_0A(256'h0000000d9ff0bb0800000014a000ba070000000d8ff2200800000014a0020779),
    .INIT_0B(256'h0000002fb2501f0000000014b000be0b0000000daff0bd0a00000014a000bc09),
    .INIT_0C(256'h0000000d1ff3243700000001a001d0c000000000200030f000000025000000e0),
    .INIT_0D(256'h00000014a04000a000000014a042247300000014a043243700000014a000d080),
    .INIT_0E(256'h00000014a04206a000000014a04206a000000014a042f01400000014a040301f),
    .INIT_0F(256'h000000062b01d07b00000020a420307f000000022a0000b000000014a04206a0),
    .INIT_10(256'h00000000b900300300000000a80000e0000000250002f0150000002f2263e473),
    .INIT_11(256'h00000014b00206a000000014a060300300000014b00000f000000014a062f013),
    .INIT_12(256'h00000014b000df0800000014a062fe1200000014b002fd1100000014a062fc10),
    .INIT_13(256'h000000002100ba130000002500003f0100000014b002f01300000014a063645d),
    .INIT_14(256'h000000032aa2fc0c00000001b003647300000001a001cab0000000003800bb02),
    .INIT_15(256'h0000000d3ff14e0600000014a002ff0f0000000d2ff2fe0e000000033012fd0d),
    .INIT_16(256'h000000002103247300000014b081df010000000daff03f0300000014a0014f00),
    .INIT_17(256'h000000033021cab0000000032cc0bb0200000001a000ba130000000038022470),
    .INIT_18(256'h00000014a002fd110000000d3ff2fc1000000014a0003e010000000d2ff36473),
    .INIT_19(256'h000000003800b206000000002100b10500000014b080b0040000000daff2fe12),
    .INIT_1A(256'h0000000d2ff3e473000000033041ae20000000032f01ad1000000001a0018c00),
    .INIT_1B(256'h0000000daff2f40f00000014a00034010000000d3ff0b40f00000014a0020b5d),
    .INIT_1C(256'h00000000950208a300000025000208fc0000002fb272068500000014b08208f8),
    .INIT_1D(256'h0000001490e2200800000001100207790000000100c2074b0000000084001000),
    .INIT_1E(256'h00000036a770d0200000001900136189000000131000d040000000148080900f),
    .INIT_1F(256'h000000018ff0900e000000019ff3618400000036a810d0800000001d10036189),
    .INIT_20(256'h000000011023617d00000036a870d0400000000d50836180000000250000d080),
    .INIT_21(256'h0000001d10336177000000250000d010000000018ff3617a000000019ff0d020),
    .INIT_22(256'h000000018ff0901b0000000004032492000000001500d0040000003ea930900e),
    .INIT_23(256'h0000003ea8c1d0e000000014008030f00000001410e2b04e000000118012f00b),
    .INIT_24(256'h000000009500d020000000250000900d00000001104224780000000190f324a1),
    .INIT_25(256'h0000003ea9c324a10000001b9041d04900000019828090060000000084036478),
    .INIT_26(256'h00000025000206da000000018ff2071e000000019ff36478000000011021d053),
    .INIT_27(256'h00000014900206dc00000014106206e00000000381f207000000000018020782),
    .INIT_28(256'h000000149002089400000014106206da000000149002070a0000001410622478),
    .INIT_29(256'h0000001d80c2f03200000036aa9010000000001d90f208a3000000011022012b),
    .INIT_2A(256'h0000003700120779000000250002074b0000000110401000000000390002d003),
    .INIT_2B(256'h0000000b40e208a30000000b30d2012b0000000b20c2089400000020b4422008),
    .INIT_2C(256'h000000144002f0320000001430001000000000142062073f0000000ba0f01060),
    .INIT_2D(256'h00000000540207790000000327f2074b000000142080100000000014a002d003),
    .INIT_2E(256'h000000006a001f000000001450e01e000000001450e01d000000000340322008),
    .INIT_2F(256'h0000001470e01d010000001470e2ff12000000007a02fe11000000036032fd10),
    .INIT_30(256'h000000008201d0ff00000001e000b00f00000001d0020b5d000000037032fd1e),
    .INIT_31(256'h00000032b0f2f00f0000001d6030300100000032ae80b00f0000001d602324cb),
    .INIT_32(256'h00000036ace0900e0000001cd30221ab00000001a002090f00000001900208f8),
    .INIT_33(256'h000000108f02f00b00000009f080901b00000032ad5324d40000001ce400d004),
    .INIT_34(256'h00000013e00324e600000011d011d0e000000013a00030f0000000139002b04e),
    .INIT_35(256'h0000000bf310bd100000000be300b20600000001d000b10500000022aca0b004),
    .INIT_36(256'h000000129f01cd00000000108e003f0100000032adf0bf120000001cd500be11),
    .INIT_37(256'h0000002f81011d0100000022ad8324e600000011d011ef2000000013a001ee10),
    .INIT_38(256'h000000140062fe110000000b0022fd1000000003a0113f000000002f91113e00),
    .INIT_39(256'h000000250002012b00000037000208940000002fa12224bf00000004a002ff12),
    .INIT_3A(256'h00000001900010000000000b2372d1030000000be31010000000000bd30208a3),
    .INIT_3B(256'h00000032af50b01e0000001cf202200800000001f002077900000001a002074b),
    .INIT_3C(256'h00000011f010b41600000013a0001200000000129e036549000000108d01d001),
    .INIT_3D(256'h0000001cf502f9170000000b23c2f81600000001f0020a7300000022aee0b517),
    .INIT_3E(256'h00000013a0020a73000000139000b519000000108200b41800000032afe04210),
    .INIT_3F(256'h0000001cf300b41a00000001f000421000000022af72f91900000011f012f818),
    .INIT_40(256'h000000138002f91b000000139002f81a0000001180220a7300000032b060b51b),
    .INIT_41(256'h0000002f91120a730000002f8100b51d00000022aff0b41c00000011f0104210),
    .INIT_42(256'h00000004a000d20200000014006042100000000b0022f91d00000003a012f81c),
    .INIT_43(256'h0000000bd3020817000000250002f21e00000037000012020000002fa123251a),
    .INIT_44(256'h000000019001d001000000018000b0320000000b2372080f0000000be3120802),
    .INIT_45(256'h00000032b1d207390000001cf20324cb00000001f001d00200000001a00324ad),
    .INIT_46(256'h00000011f012f21e00000013a0001204000000129e02258a000000108d005020),
    .INIT_47(256'h0000001df002f01400000003ff00b1170000000bf390b01600000022b1620c13),
    .INIT_48(256'h0000001df02346850000000b23c1f1ff00000001f001d0ff00000032b2a2f115),
    .INIT_49(256'h00000013a002f115000000139002f014000000108200b11900000032b2a0b018),
    .INIT_4A(256'h0000000b2380b01a00000001f003468500000022b231f1ff00000011f011d0ff),
    .INIT_4B(256'h000000139001d0ff000000108202f11500000032b332f0140000001cf500b11b),
    .INIT_4C(256'h00000001f000b11d00000022b2c0b01c00000011f013468500000013a001f1ff),
    .INIT_4D(256'h000000139001f1ff000000118011d0ff00000032b3b2f1150000001cf302f014),
    .INIT_4E(256'h0000002f8103653d00000022b341d00000000011f010b0320000001380034685),
    .INIT_4F(256'h000000140062083e0000000b0022080200000003a01208170000002f911208fc),
    .INIT_50(256'h00000025000324ad000000370001d0010000002fa120b03200000004a002080f),
    .INIT_51(256'h0000002f504030df000000096082073900000009508324cb00000020b561d002),
    .INIT_52(256'h0000002f530206fe0000000960836556000000095081d0080000002f6052258a),
    .INIT_53(256'h0000002f537207e700000009608206da00000009508206fe0000002f6312071c),
    .INIT_54(256'h0000002f53c2073900000009608324ad000000095081d0010000002f6380b032),
    .INIT_55(256'h0000000160736563000000015f01d010000000250002258a0000002f60605020),
    .INIT_56(256'h0000002d10b206da0000002d60a207280000002d5092072200000001100206fa),
    .INIT_57(256'h0000000b810324ad00000020b441d001000000370010b03200000025000207e7),
    .INIT_58(256'h0000002f9351d0200000002f8342258a0000000ba12050200000000b91120739),
    .INIT_59(256'h0000000b330207280000000bd372072200000001200206fa0000002fa3636570),
    .INIT_5A(256'h0000001ba001d0010000001a9400b03200000018830207e70000000b431206da),
    .INIT_5B(256'h0000002f9352258a0000002f834030df00000011201207390000003ab74324ad),
    .INIT_5C(256'h00000022b692072200000032ba6206fa0000001c2d03657d0000002fa361d040),
    .INIT_5D(256'h0000002f20f0b0320000000ba36207e70000000b935206da0000000b83420728),
    .INIT_5E(256'h0000001d401030df000000094082073900000001300324ad000000012001d001),
    .INIT_5F(256'h0000001ba002071c0000001b90036017000000188401d08000000032c0c2258a),
    .INIT_60(256'h0000002f834207e700000013300206da00000011201207120000003ab8720716),
    .INIT_61(256'h0000000b8342073900000022b7a324ad0000002fa361d0010000002f9350b032),
    .INIT_62(256'h0000002f20d010080000002f30e2073f0000000ba362258a0000000b935030df),
    .INIT_63(256'h000000144061d0040000000b50d0b01e0000000b40c220080000002f80c2074b),
    .INIT_64(256'h0000000b50d325ed0000002f40c0d00400000014408090020000001450836602),
    .INIT_65(256'h0000002f50d0bf05000000145080be0400000014608206740000000b60e2064e),
    .INIT_66(256'h0000001460801f0900000014608325a00000000b70f1ff320000000b60e1dedb),
    .INIT_67(256'h00000001700225a40000002f70e0120b0000000377f011bb0000001470001ed0),
    .INIT_68(256'h0000002f70f0120c000000047000112b0000001400601e400000000b00201f0a),
    .INIT_69(256'h000000034f02de090000000b4392df0a0000002500009d070000003700020626),
    .INIT_6A(256'h000000012001cf200000000b43c365ae00000032bdd1ce100000001d4002dd08),
    .INIT_6B(256'h0000003abb713f000000001ba0011e010000001b900225b100000018840365ae),
    .INIT_6C(256'h0000002fa362f0140000002f9350b1170000002f8340b01600000011201225a4),
    .INIT_6D(256'h0000000b834325bd00000022bac1f1ff00000032bdd1d0ff0000001d2022f115),
    .INIT_6E(256'h0000000b43c142000000002f20f0d0ff0000000ba36012000000000b9352062e),
    .INIT_6F(256'h0000001ba002f0140000001b9000b119000000188400b018000000194022f220),
    .INIT_70(256'h0000000ba36325c90000000b9351f1ff0000000b8341d0ff0000003ec0c2f115),
    .INIT_71(256'h0000001490e14200000000033010d0ff00000000380012000000000b20f2062e),
    .INIT_72(256'h000000143082f014000000148080b11b000000143060b01a000000148082f221),
    .INIT_73(256'h00000014808325d5000000149081f1ff000000148061d0ff0000002f30c2f115),
    .INIT_74(256'h0000001420614200000000142000d0ff00000014908012000000002f80d2062e),
    .INIT_75(256'h0000000b00201200000000013010b11d0000002f20e0b01c0000001420e2f222),
    .INIT_76(256'h000000370001f1ff0000002f30f1d0ff000000043002f115000000140062f014),
    .INIT_77(256'h000000188400d0ff00000001200012000000000b4382062e00000025000325e2),
    .INIT_78(256'h00000011201208570000003abe82080a0000001ba002f2230000001b90014200),
    .INIT_79(256'h00000022bdf040100000002fa360b1210000002f9350b0200000002f8342080f),
    .INIT_7A(256'h0000002f20f040100000000ba360b1230000000b935040100000000b8340b122),
    .INIT_7B(256'h0000001b900225f2000000188400504000000019402207390000000b438325f0),
    .INIT_7C(256'h0000000b9350b00e0000000b8342073f0000003ec0c030bf0000001ba0020739),
    .INIT_7D(256'h00000014808365fe0000000b300190010000000b20f0b01f0000000ba362f03b),
    .INIT_7E(256'h000000149082b80f000000148062b40f0000002f30c2b20f00000014308208a3),
    .INIT_7F(256'h0000001420001082000000149082f01f0000002f80d226230000001480801002),
    .INITP_00(256'h02b91f291fa83c0e3c083c8bba14231a901191288aa69a2799243800af1715a7),
    .INITP_01(256'h0a9a3e0c0c0c84931a19829f9ba7a1af17a6a10e228b83971494a6b385ba0a37),
    .INITP_02(256'h94aaa12629253e9f300d01141881a2a6bebd3b8e2a0cad873300a79f1a2db98e),
    .INITP_03(256'h8021a32fa03f9f391e1337153ca19c3b3b8d3d85101ea338bca6ac2f8ea11205),
    .INITP_04(256'h1e3dac933895a69e8b1d0601a3279c3a851ab7a60c3c89902e3882b91ea3b83d),
    .INITP_05(256'h38bc9202b31c1f28309a2982b6973eb41c2885b32cb30a88b92c0c0e02bc1e22),
    .INITP_06(256'h8c15253b008eb539349a1b11103e23ad999ba33b1e87a9279e0d3f8e3f130225),
    .INITP_07(256'hbd301f1a20ba0726110d251f03ba119630b0b43430128b82b324a42d88b31d26),
    .INITP_08(256'h1399b93a863c129c17a8a33c24931c9a8bb6b8bc33163e99a705978101acb797),
    .INITP_09(256'h043d98a21dbd809fb936053531278f3ea7841602023ea3943039068d0d992581),
    .INITP_0A(256'h84b6a9342d991d94b8afaaaaba8890afac0b8029319414af320d8db5bb27b52a),
    .INITP_0B(256'h1f848fa538a9398596373d0808a41faaaa932e818a9fb001b50d13282d932e38),
    .INITP_0C(256'h83059cac95880aa4311b06a7a711381ba3a102968a22a9af021a22b00db9a50a),
    .INITP_0D(256'h941f1c8b8c943d3f03018e263c328534901b8180038686bab81db63e9f9f8cb3),
    .INITP_0E(256'h169f843ab9a1b89d222802aa2d3686052202253000281da91182b919b2bf98b8),
    .INITP_0F(256'hbd83142e0f28ac9e3db01b34370127908c0b048899b4ba08a534bc1ab6a11907),
