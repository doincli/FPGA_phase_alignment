    .INIT_00(256'h0142083261d200200143081d0022ff000013032200801f000142062076128000),
    .INIT_01(256'h0140063261d2074b00b0021d010010010013013261d2004902f20e1d00820033),
    .INIT_02(256'h025000050401d002037000207393205d02f30f3660f1d0010043001d0202073c),
    .INIT_03(256'h02f20e1d0401d01002f20d226233226302f20c010021d0000012ff2073f32143),
    .INIT_04(256'h0013002073f1d008025000030bf324ef037000207391d00402f20f366163242a),
    .INIT_05(256'h02f0163601701060020c301d0803222a00b117226231d08200b016010023258e),
    .INIT_06(256'h00b01801002207080013012073f2074b02f220030bf0109f02f117207392073f),
    .INIT_07(256'h02f1192073922ffd02f018208a3206da020c302012b2072000b1192262320710),
    .INIT_08(256'h00b11b2074b0b00000b01a010003202f0013022073f0d08002f2210504009002),
    .INIT_09(256'h02f2220d080011ff02f11b0900d010ff02f01a220083602f020c30207790d001),
    .INIT_0A(256'h020c300d0401b20000b11d0900d1b10000b01c2500019001001303366260121f),
    .INIT_0B(256'h025000015090900102f223014d02f00002f11d250000100102f01c3662a3e029),
    .INIT_0C(256'h0310001ff322b00001f1ff1dedb2500001d0ff0bf053202f0012000be040d040),
    .INIT_0D(256'h0140060150a09001014006014402be0f014006226382bf7e014006326362b00c),
    .INIT_0E(256'h01400e0d0100d0200141000b0140900d0140060b2152d001014100013000300f),
    .INIT_0F(256'h00b22414200090060100300d0082203a01400e143000900601400e142003603f),
    .INIT_10(256'h022ffd1900136046022ffd011010d080022ffd030070900d0250001430009006),
    .INIT_11(256'h022ffd1024009007022ffd2264309007022ffd1410622041022ffd3a64709007),
    .INIT_12(256'h022ffd0900820712022ffd2d20920702022ffd2d30a2071e022ffd1235025000),
    .INIT_13(256'h022ffd0bb1320720022ffd01a0020710022ffd2500020722022ffd02010206de),
    .INIT_14(256'h022ffd09d1d20724022ffd09c1c206de022ffd14b06206fa022ffd14b062071c),
    .INIT_15(256'h022ffd10cb0206da022ffd10ba0206e2022ffd09f1f206de022ffd09e1e206e4),
    .INIT_16(256'h022ffd01a043e05a022ffd13f0019001022ffd13e0001019022ffd13d0025000),
    .INIT_17(256'h022ffd09c07200da022ffd20626200f4022ffd20678200ec022ffd01b0025000),
    .INIT_18(256'h022ffd09e0720894022ffd2062632060022ffd09d070d001022ffd206260900d),
    .INIT_19(256'h022ffd01b01208b5022ffd01aeb208d2022ffd09f0701101022ffd2062601080),
    .INIT_1A(256'h022ffd0360101000022ffd0b61236063022ffd0b5111dc93022ffd0b410208e2),
    .INIT_1B(256'h022ffd13f002f002022ffd12e6001000022ffd12d502f001022ffd10c4005001),
    .INIT_1C(256'h022ffd250001d102022ffd3e66c0311e022ffd1bb00001e0022ffd19a0120b44),
    .INIT_1D(256'h022ffd250001d104022ffd2067832080022ffd01b011d110022ffd01aec3207e),
    .INIT_1E(256'h022ffd2de071d116022ffd2062a32087022ffd2df071d112022ffd2062a32085),
    .INIT_1F(256'h022ffd2dc073209f022ffd2062a01200022ffd2dd0722017022ffd2062a3208b),
    .INIT_20(256'h022ffd2da073209f022ffd2062a1d190022ffd2db0701220022ffd2062a001d0),
    .INIT_21(256'h022ffd01300001d0022ffd015003209f022ffd0146c01203022ffd250002208b),
    .INIT_22(256'h022ffd1420001000022ffd0d0103209f022ffd0b0141d190022ffd0b21501204),
    .INIT_23(256'h022ffd1430014000022ffd142000dd40022ffd0d00836092022ffd143000dd10),
    .INIT_24(256'h022ffd3a6961d110022ffd190012f002022ffd0110114000022ffd030070dd20),
    .INIT_25(256'h022ffd123501d116022ffd102403209b022ffd226921d112022ffd1410632099),
    .INIT_26(256'h022ffd0601001223022ffd090083209f022ffd2d20901222022ffd2d30a3209d),
    .INIT_27(256'h022ffd250002f239022ffd2d0083209f022ffd2d20901226022ffd2d30a3209f),
    .INIT_28(256'h022ffd14d0009002022ffd14c002f03a022ffd14b0001000022ffd14a06200d6),
    .INIT_29(256'h022ffd110b9200e6022ffd250002f024022ffd14f0001001022ffd14e000d004),
    .INIT_2A(256'h022ffd19011208a3022ffd390002089d022ffd190e9208a0022ffd39000200ff),
    .INIT_2B(256'h022ffd190f62090b022ffd390002b02e022ffd110072090b022ffd3e6b12b02e),
    .INIT_2C(256'h022ffd00c002011d022ffd25000200e0022ffd1100a200d6022ffd2500020894),
    .INIT_2D(256'h022ffd206bb0300f022ffd2072e09001022ffd206c52b04e022ffd206bb200d6),
    .INIT_2E(256'h022ffd011000d002022ffd2500009002022ffd2072e320cb022ffd206c51d001),
    .INIT_2F(256'h022ffd141002b40f022ffd14c062b20f022ffd14100208a3022ffd14c06320c5),
    .INIT_30(256'h022ffd1410020779022ffd14c062074b022ffd1410001002022ffd14c062b80f),
    .INIT_31(256'h022ffd1110701000022ffd3a6c8208a3022ffd1d10a2012b022ffd2500022008),
    .INIT_32(256'h022ffd20731208a3022ffd01a0022008022ffd2500020779022ffd111302074b),
    .INIT_33(256'h022ffd0110401001022ffd390002b80f022ffd206a72b40f022ffd090062b20f),
    .INIT_34(256'h022ffd04a00206e0022ffd366d020700022ffd1910120767022ffd206a02f032),
    .INIT_35(256'h022ffd192012070e022ffd2072e20716022ffd206c522478022ffd00100206dc),
    .INIT_36(256'h022ffd2272e206fe022ffd0110d2070a022ffd2500025000022ffd366cb206da),
    .INIT_37(256'h022ffd2272e25000022ffd0115f206dc022ffd2272e20718022ffd01120206fa),
    .INIT_38(256'h022ffd2272e20720022ffd011312070a022ffd2272e20714022ffd0113e2070a),
    .INIT_39(256'h022ffd2272e20700022ffd011302071c022ffd2272e25000022ffd01133206dc),
    .INIT_3A(256'h022ffd2272e25000022ffd01132206dc022ffd2272e2070e022ffd01131206fc),
    .INIT_3B(256'h022ffd2272e09001022ffd01134206dc022ffd2272e2071e022ffd0113320704),
    .INIT_3C(256'h022ffd2272e25000022ffd01136206da022ffd2272e206b3022ffd011350300f),
    .INIT_3D(256'h022ffd2272e09002022ffd01138206dc022ffd2272e20704022ffd01137206fa),
    .INIT_3E(256'h022ffd2272e1400e022ffd011411400e022ffd2272e1400e022ffd0113903008),
    .INIT_3F(256'h022ffd2272e010c0022ffd0114325000022ffd2272e206da022ffd01142206b3),
    .INIT_40(256'h022ffd2272e01e00022ffd0114501f00022ffd2272e208d2022ffd0114401100),
    .INIT_41(256'h022ffd2272e010a0022ffd01147208ec022ffd2272e01c00022ffd0114601d01),
    .INIT_42(256'h022ffd2272e01e00022ffd0114901f00022ffd2272e208d2022ffd0114801100),
    .INIT_43(256'h022ffd2272e010c0022ffd0114b208ec022ffd2272e01c00022ffd0114a01d00),
    .INIT_44(256'h022ffd2272e03f81022ffd0114d208e9022ffd2272e208d2022ffd0114c01101),
    .INIT_45(256'h022ffd2272e05f00022ffd0114f03c3f022ffd2272e03d7c022ffd0114e03e3c),
    .INIT_46(256'h022ffd2272e208ec022ffd0115105c00022ffd2272e05d03022ffd0115005e40),
    .INIT_47(256'h022ffd2272e208d2022ffd0115301101022ffd2272e010c0022ffd0115225000),
    .INIT_48(256'h022ffd2272e03dfd022ffd0115503e7f022ffd2272e03fff022ffd01154208e9),
    .INIT_49(256'h022ffd2272e05d00022ffd0115705e80022ffd2272e05f00022ffd0115603cff),
    .INIT_4A(256'h022ffd2272e010c0022ffd0115925000022ffd2272e208ec022ffd0115805c00),
    .INIT_4B(256'h022ffd2d10603fff022ffd20735208e9022ffd2272e208d2022ffd0115a01101),
    .INIT_4C(256'h022ffd36731208ec022ffd0d02003cff022ffd0900d03dfe022ffd2500003eff),
    .INIT_4D(256'h022ffd36735208d2022ffd0d01001101022ffd0900d010c0022ffd2500025000),
    .INIT_4E(256'h022ffd2500003dfe022ffd0306003eff022ffd0900003fff022ffd25000208e9),
    .INIT_4F(256'h022ffd0010005d01022ffd2500005e00022ffd0309f05f00022ffd0900003cff),
    .INIT_50(256'h022ffd2d10001000022ffd0410025000022ffd2073c208ec022ffd0316005c00),
    .INIT_51(256'h022ffd207390d040022ffd206dc0900f022ffd206fe2f01e022ffd207042f032),
    .INIT_52(256'h022ffd001000d080022ffd2500036189022ffd206da0d020022ffd206b336189),
    .INIT_53(256'h022ffd2d10036180022ffd041000d080022ffd207390900e022ffd0319f36184),
    .INIT_54(256'h022ffd0b0323617a022ffd206dc0d020022ffd206fe3617d022ffd2071e0d040),
    .INIT_55(256'h022ffd206b30d004022ffd2073c0900e022ffd3277536177022ffd1d0010d010),
    .INIT_56(256'h022ffd206fe2b04e022ffd2071e2f00b022ffd250000901b022ffd206da32160),
    .INIT_57(256'h022ffd206da2216e022ffd206b33616d022ffd010021d0e0022ffd206dc030f0),
    .INIT_58(256'h022ffd2073909006022ffd0319f3616d022ffd001000d020022ffd250000900d),
    .INIT_59(256'h022ffd010001d053022ffd250002216e022ffd2d10036167022ffd041001d049),
    .INIT_5A(256'h022ffd2071e20782022ffd2d103206da022ffd0b1322071e022ffd207613616d),
    .INIT_5B(256'h022ffd1d001206da022ffd0b0322070a022ffd206dc22008022ffd206fe20779),
    .INIT_5C(256'h022ffd206da01000022ffd206b3208a3022ffd010402012b022ffd3277520894),
    .INIT_5D(256'h022ffd206da2b10e022ffd206b322008022ffd0102020779022ffd250002074b),
    .INIT_5E(256'h022ffd3278001040022ffd1d0002b20e022ffd2073c22187022ffd2500001080),
    .INIT_5F(256'h022ffd2500022187022ffd206dc01020022ffd206e02b40e022ffd2071622187),
    .INIT_60(256'h022ffd2071422187022ffd2071e01010022ffd2277d2b80e022ffd2070a20894),
    .INIT_61(256'h022ffd206da2f01e022ffd206b401008022ffd0bc022b80f022ffd206dc20894),
    .INIT_62(256'h022ffd2070a2b20f022ffd2071c2b40f022ffd2074420894022ffd2075022200),
    .INIT_63(256'h022ffd206da19801022ffd206b40982f022ffd0bc3a2f01e022ffd206dc01001),
    .INIT_64(256'h022ffd206dc208d2022ffd2070401102022ffd20712010a0022ffd250000b203),
    .INIT_65(256'h022ffd206b42fc0c022ffd0bc0603f03022ffd206e6208e2022ffd206e6208b5),
    .INIT_66(256'h022ffd206b40bc0c022ffd0bc042ff0f022ffd206b42fe0e022ffd0bc052fd0d),
    .INIT_67(256'h022ffd206fc01020022ffd207200bf0f022ffd207e70be0e022ffd206da0bd0d),
    .INIT_68(256'h022ffd3a7a60b001022ffd0d504208ec022ffd09502208d2022ffd206dc01100),
    .INIT_69(256'h022ffd09d1d221ab022ffd09c1c22017022ffd227bd361a8022ffd207f90d001),
    .INIT_6A(256'h022ffd14b060b016022ffd0bb022090f022ffd09f1f208c1022ffd09e1e208a9),
    .INIT_6B(256'h022ffd13e000b018022ffd13d001f000022ffd10cb00b017022ffd14b061d000),
    .INIT_6C(256'h022ffd2fd350b01a022ffd2fe361f000022ffd2ff3b0b019022ffd13f001f000),
    .INIT_6D(256'h022ffd0bc360b01c022ffd206b41f000022ffd0bc3b0b01b022ffd2fc341f000),
    .INIT_6E(256'h022ffd0bc34361c7022ffd206b41f000022ffd0bc350b01d022ffd206b41f000),
    .INIT_6F(256'h022ffd206fc0b03a022ffd206fe324cb022ffd206da1d002022ffd206b40b032),
    .INIT_70(256'h022ffd207f90b032022ffd3a7c5208a3022ffd0d5042f03a022ffd206dc11001),
    .INIT_71(256'h022ffd0be360b001022ffd0bd3522008022ffd0bc3432478022ffd227db1d001),
    .INIT_72(256'h022ffd20678321fd022ffd01b001d800022ffd01a04308f8022ffd0bf3b0d001),
    .INIT_73(256'h022ffd09e072f035022ffd206260b017022ffd09f072f034022ffd206260b016),
    .INIT_74(256'h022ffd09c072f03b022ffd206260b019022ffd09d072f036022ffd206260b018),
    .INIT_75(256'h022ffd00ce02f03d022ffd206b40b01b022ffd00cd02f03c022ffd206b40b01a),
    .INIT_76(256'h022ffd206da2f03f022ffd206b40b01d022ffd00cf02f03e022ffd206b40b01c),
    .INIT_77(256'h022ffd206e62090f022ffd206dc208c1022ffd20710208a9022ffd206fe208ef),
    .INIT_78(256'h022ffd11c010b017022ffd14c001c010022ffd0d5040b134022ffd01c000b016),
    .INIT_79(256'h022ffd207200b136022ffd250000b018022ffd206da1e010022ffd206b40b135),
    .INIT_7A(256'h022ffd2b03c1e010022ffd2b80c0b13b022ffd206dc0b019022ffd2071e1e010),
    .INIT_7B(256'h022ffd09c0c0b01b022ffd2b02c1e010022ffd206b40b13c022ffd09c0c0b01a),
    .INIT_7C(256'h022ffd206b40b13e022ffd09c0c0b01c022ffd2b01c1e010022ffd206b40b13d),
    .INIT_7D(256'h022ffd206da1e010022ffd206b40b13f022ffd09c0c0b01d022ffd2b00c1e010),
    .INIT_7E(256'h022ffd20728321fd022ffd207281d800022ffd2072819801022ffd250003620f),
    .INIT_7F(256'h022ffd207282f01f022ffd2072801004022ffd2072820aab022ffd20728221dc),
    .INITP_00(256'h4b68d82918057578617c042f397ccf6aecd14786685ed7bbb989a8ce3ea13d93),
    .INITP_01(256'h2604b09592971d93a0b408297faca785e55e5e76cc88b92663eb66fc37b0144b),
    .INITP_02(256'hd179d24ef3eb45ccc8f052ea66546d6ed36e6ff3deec46f370fbf366ebd8ce46),
    .INITP_03(256'hdff16172e9f34c76f5d744fff64af6efeb51d155dff966c9497151f2ebff7969),
    .INITP_04(256'h65dc67c0d6d9e145e0e17fec67f7c5c15ef466556df373dafa68fe725e607b6e),
    .INITP_05(256'h73557ecfcb7946f74d567dd1cbe149fef05e42c07dd26447e8e0ce69794e68c4),
    .INITP_06(256'h6bfb6f526c5feadb5ec3756369d8dcd850c65f59ca7fec66f9c5e2f8efce6fca),
    .INITP_07(256'hefec60f87c607cddf8d867516bc165dcfe596cc06bdee5d5e1cf6bc46b5fee5f),
    .INITP_08(256'h77ffef687060e97fe1e7e1f569e87761ef6a767b78f477fe6eeb76797875777f),
    .INITP_09(256'h6c6df1c869facbf477ffdaea6cfedde96a5f7778ef7470e7ef65e179ee7a65f1),
    .INITP_0A(256'he35eed6de04574f143d4f15667f1edcbf54cd2c8657876d54968f65ae042dd53),
    .INITP_0B(256'hfe70e0cb6fdfd265e555f66a7dd0cef7567feb7bc169537bff777859d54163fe),
    .INITP_0C(256'h6f46566a40eec87f43e26163e551c6e76c506279db436fe2f5de71ed50c8d2d4),
    .INITP_0D(256'h62776f596e5d675d655d7e71c14e79efc04bcf78634a4cf3ffc54dc253ed44f7),
    .INITP_0E(256'h636a4d60fc54c8d7505752d45f757ef6ff715ff2d04b73754ad870f8407d716f),
    .INITP_0F(256'h4cc1dad3cc4156f4e256c95cd54ac2d3ca435049ddecf1ded161e2d451467b63),
