    .INIT_00(256'h022ffd1d0001d002022ffd0b0320b032022ffd250002f013022ffd207280b002),
    .INIT_01(256'h022ffd2071c0b032022ffd207162078a022ffd206fe206da022ffd3680932206),
    .INIT_02(256'h022ffd20710324ef022ffd206fe1d002022ffd25000324ef022ffd206da1d001),
    .INIT_03(256'h022ffd0b0320b03a022ffd2500022008022ffd206da2074b022ffd206fa01004),
    .INIT_04(256'h022ffd207141d000022ffd207020b016022ffd368162f03a022ffd1d00011001),
    .INIT_05(256'h022ffd207021f000022ffd250000b018022ffd206da1f000022ffd207000b017),
    .INIT_06(256'h022ffd207e71f000022ffd206da0b01a022ffd206fe1f000022ffd206fe0b019),
    .INIT_07(256'h022ffd0b1131f000022ffd206dc0b01c022ffd206fa1f000022ffd207180b01b),
    .INIT_08(256'h022ffd00c00208a3022ffd0401036017022ffd0b00f1f000022ffd141060b01d),
    .INIT_09(256'h022ffd2072e1d002022ffd206c532478022ffd206bb1d001022ffd206bb0b032),
    .INIT_0A(256'h022ffd206b32f01e022ffd0b00d01001022ffd206b322008022ffd0b00e324cb),
    .INIT_0B(256'h022ffd2071011d01022ffd206da0bf12022ffd206b30be11022ffd0b00c0bd10),
    .INIT_0C(256'h022ffd0b1132fe11022ffd206e62fd10022ffd206dc13f00022ffd206fa13e00),
    .INIT_0D(256'h022ffd206b30b00f022ffd0401020b5d022ffd0b0122ff12022ffd1410603f01),
    .INIT_0E(256'h022ffd206b30307e022ffd0b0100b03b022ffd206b32f00f022ffd0b01103001),
    .INIT_0F(256'h022ffd1dcff3625b022ffd0bc171c0e0022ffd2500003e7e022ffd206da0be0e),
    .INIT_10(256'h022ffd348821d000022ffd1dcff0b016022ffd0bc162090f022ffd3487c208f8),
    .INIT_11(256'h022ffd0bc181f000022ffd3487c0b018022ffd1dcff1f000022ffd0bc190b017),
    .INIT_12(256'h022ffd1dcff1f000022ffd0bc1b0b01a022ffd348821f000022ffd1dcff0b019),
    .INIT_13(256'h022ffd348821f000022ffd1dcff0b01c022ffd0bc1a1f000022ffd3487c0b01b),
    .INIT_14(256'h022ffd0bc1c2225b022ffd3487c36254022ffd1dcff1f000022ffd0bc1d0b01d),
    .INIT_15(256'h022ffd0bd202078a022ffd25000206da022ffd3488220779022ffd1dcff2075a),
    .INIT_16(256'h022ffd2087c208a3022ffd0bc1722008022ffd328602074b022ffd1dd0001004),
    .INIT_17(256'h022ffd2088e01002022ffd0bc202b80f022ffd208882b40f022ffd0bc162b20f),
    .INIT_18(256'h022ffd0bc1901000022ffd3286922008022ffd1dd0020779022ffd0bd212074b),
    .INIT_19(256'h022ffd0bc2132294022ffd208880d004022ffd0bc180900e022ffd2087c2f032),
    .INIT_1A(256'h022ffd328722f008022ffd1dd0009018022ffd0bd222f007022ffd2088e09017),
    .INIT_1B(256'h022ffd208882f00a022ffd0bc1a0901a022ffd2087c2f009022ffd0bc1b09019),
    .INIT_1C(256'h022ffd1dd00030f0022ffd0bd232b04e022ffd2088e2f00b022ffd0bc220901b),
    .INIT_1D(256'h022ffd0bc1c0d002022ffd2087c09002022ffd0bc1d3627a022ffd3287b1d0a0),
    .INIT_1E(256'h022ffd250003627d022ffd2088e1d0e0022ffd0bc23223ed022ffd20888323ec),
    .INIT_1F(256'h022ffd206b40bc07022ffd206dc36287022ffd207001d0b0022ffd20726223ec),
    .INIT_20(256'h022ffd20720206dc022ffd206fc2071c022ffd250002dc01022ffd206dc03c0f),
    .INIT_21(256'h022ffd250001d0d0022ffd206da22003022ffd206b4206da022ffd206dc206b4),
    .INIT_22(256'h022ffd206b41d0f0022ffd206dc22409022ffd2072020722022ffd206fc3628b),
    .INIT_23(256'h022ffd207241d0c0022ffd20710223f9022ffd2500020700022ffd206dc3628f),
    .INIT_24(256'h022ffd25000223ea022ffd206da32412022ffd206b40d080022ffd206dc32412),
    .INIT_25(256'h022ffd2b08e09006022ffd2b1bb363ec022ffd2b00a0d020022ffd2b0090900d),
    .INIT_26(256'h022ffd200590d002022ffd208ac09002022ffd01c003629e022ffd209071d04f),
    .INIT_27(256'h022ffd25000362a5022ffd208ac1d053022ffd01c10223ed022ffd25000323ec),
    .INIT_28(256'h022ffd01c0d20791022ffd2500020782022ffd208ac206da022ffd01c072071e),
    .INIT_29(256'h022ffd208ac2071c022ffd01c01362bc022ffd250001d052022ffd208ac223eb),
    .INIT_2A(256'h022ffd25000363ea022ffd208ac1d020022ffd01c0409006022ffd2500020731),
    .INIT_2B(256'h022ffd208db1d030022ffd01f0009006022ffd01e0020731022ffd01d00206dc),
    .INIT_2C(256'h022ffd208bb09006022ffd208d220731022ffd01100206e6022ffd01080363ea),
    .INIT_2D(256'h022ffd2b63b00100022ffd2b00a2d001022ffd2b3893a3ea022ffd25000206a7),
    .INIT_2E(256'h022ffd2b1c922003022ffd25000206da022ffd209072072e022ffd2b08e206c5),
    .INIT_2F(256'h022ffd2090722409022ffd2b08e20722022ffd2b37b362c0022ffd2b00a1d055),
    .INIT_30(256'h022ffd2b0bb223f9022ffd2b72a20700022ffd2b649362c4022ffd250001d044),
    .INIT_31(256'h022ffd2b64920731022ffd2500020714022ffd20907362d5022ffd2b08e1d04e),
    .INIT_32(256'h022ffd20907206dc022ffd2b08e363ea022ffd2b57b1d020022ffd2b20a09006),
    .INIT_33(256'h022ffd2b08e2fa07022ffd2b63b3a3ea022ffd2b20a206ca022ffd2b6c90120a),
    .INIT_34(256'h022ffd2b4192fe0b022ffd2b00a2fd0a022ffd250002fc09022ffd209072fb08),
    .INIT_35(256'h022ffd2b25920720022ffd2b00a36328022ffd2d1081d054022ffd2d0082241e),
    .INIT_36(256'h022ffd2b00a363ea022ffd250001d020022ffd2d10809006022ffd2d00820731),
    .INIT_37(256'h022ffd2de083a3ea022ffd2dd08206ca022ffd2dc080120a022ffd2b289206dc),
    .INIT_38(256'h022ffd2b28932306022ffd2b00a1dec0022ffd250002fb3f022ffd2df082fa3e),
    .INIT_39(256'h022ffd09f08206a0022ffd09e08223ea022ffd09d08322e7022ffd09c080de80),
    .INIT_3A(256'h022ffd2500018fa0022ffd208e20ba02022ffd208b5206a0022ffd25000206a0),
    .INIT_3B(256'h022ffd010202fd0d022ffd250002fc0c022ffd208bb206a0022ffd208db363ea),
    .INIT_3C(256'h022ffd0be0e206da022ffd0bf0f20aab022ffd208d22ff0f022ffd011002fe0e),
    .INIT_3D(256'h022ffd25000206fe022ffd208ec0bf12022ffd0bc0c0be11022ffd0bd0d0bd10),
    .INIT_3E(256'h022ffd25000206b4022ffd208c100ce0022ffd208a9206b4022ffd208ef00cf0),
    .INIT_3F(256'h022ffd01080206bb022ffd208ef0bc3f022ffd25000206b4022ffd208fe00cd0),
    .INIT_40(256'h022ffd208bb0bc3e022ffd208b52072e022ffd208d2206c5022ffd01101206bb),
    .INIT_41(256'h022ffd0900e206a0022ffd25000206a0022ffd208c7223ea022ffd208a6206b4),
    .INIT_42(256'h022ffd0900e363ea022ffd2500018ea0022ffd369070ba02022ffd0d008206a0),
    .INIT_43(256'h022ffd370012fe12022ffd250002fd11022ffd3290b2fc10022ffd0d002206a0),
    .INIT_44(256'h022ffd2f1180be0d022ffd2f1170bf0c022ffd2f116206da022ffd0110020b5d),
    .INIT_45(256'h022ffd2f11c206bb022ffd2f11b206bb022ffd2f11a0bc0f022ffd2f1190bd0e),
    .INIT_46(256'h022ffd2b00a206b4022ffd2b6c900cd0022ffd010842072e022ffd2f11d206c5),
    .INIT_47(256'h022ffd2092a206b4022ffd2092500cf0022ffd11001206b4022ffd2b00b00ce0),
    .INIT_48(256'h022ffd37000206c5022ffd3691d206bb022ffd1d0ff206bb022ffd209840bc3f),
    .INIT_49(256'h022ffd09e08223ea022ffd09d08206b4022ffd09c080bc3e022ffd250002072e),
    .INIT_4A(256'h022ffd329400d004022ffd1d0c109002022ffd2500036346022ffd09f081d058),
    .INIT_4B(256'h022ffd2097309006022ffd001f020731022ffd3295520728022ffd1d0c23e346),
    .INIT_4C(256'h022ffd2097301208022ffd001d0206dc022ffd20973363ea022ffd001e01d020),
    .INIT_4D(256'h022ffd2f1282fa34022ffd01100206da022ffd209733a3ea022ffd001c0206ca),
    .INIT_4E(256'h022ffd2f1290bc34022ffd2f12e2fd3b022ffd2f12c2fc36022ffd2f12a2fb35),
    .INIT_4F(256'h022ffd2500001a01022ffd2f12f0bf3b022ffd2f12d0be36022ffd2f12b0bd35),
    .INIT_50(256'h022ffd2097309c07022ffd001e020626022ffd2097320678022ffd001f001b00),
    .INIT_51(256'h022ffd209733638e022ffd001c01d051022ffd20973223ea022ffd001d0206b4),
    .INIT_52(256'h022ffd2f42e1d020022ffd2f52c09006022ffd2f62a20731022ffd2f7282071a),
    .INIT_53(256'h022ffd01700206ca022ffd016000120a022ffd01500206dc022ffd01400363ea),
    .INIT_54(256'h022ffd2f42f0de80022ffd2f52d32362022ffd2f62b1dec0022ffd2f7293a3ea),
    .INIT_55(256'h022ffd001e0206a0022ffd20973206a0022ffd001f0223ea022ffd2293f32356),
    .INIT_56(256'h022ffd001c0363ea022ffd2097318fa0022ffd001d00ba02022ffd20973206a0),
    .INIT_57(256'h022ffd2f1292fe0e022ffd0310f2fd0d022ffd001702fc0c022ffd20973206a0),
    .INIT_58(256'h022ffd2f12b206a0022ffd0310f206a0022ffd0016022378022ffd037f02ff0f),
    .INIT_59(256'h022ffd2f12d363ea022ffd0310f18ea0022ffd001500ba02022ffd036f0206a0),
    .INIT_5A(256'h022ffd2f12f2fe12022ffd0310f2fd11022ffd001402fc10022ffd035f0206a0),
    .INIT_5B(256'h022ffd2f12a18c00022ffd2f1280b206022ffd011000b105022ffd034f00b004),
    .INIT_5C(256'h022ffd1410020b5d022ffd2293f3e3ea022ffd2f12e1ae20022ffd2f12c1ad10),
    .INIT_5D(256'h022ffd1410022378022ffd145002f40f022ffd1410003401022ffd144000b40f),
    .INIT_5E(256'h022ffd141002b00a022ffd14700206da022ffd14100208f8022ffd1460020894),
    .INIT_5F(256'h022ffd1410009e08022ffd1450009f08022ffd141000127b022ffd144002b6c9),
    .INIT_60(256'h022ffd2500000cd0022ffd14700206b4022ffd1410009c08022ffd1460009d08),
    .INIT_61(256'h022ffd20a2500cf0022ffd0b929206b4022ffd0b82800ce0022ffd00170206b4),
    .INIT_62(256'h022ffd0ba253637e022ffd01b0019201022ffd20a4f206da022ffd20a31206b4),
    .INIT_63(256'h022ffd14a00363ec022ffd0ba261d050022ffd14b00223eb022ffd14a0e208a3),
    .INIT_64(256'h022ffd14a001d020022ffd14b0009006022ffd14a0020731022ffd14b0020718),
    .INIT_65(256'h022ffd2f217206ca022ffd062b001202022ffd0b217206dc022ffd14b00363ea),
    .INIT_66(256'h022ffd14b00206a0022ffd14a00206a0022ffd14b00206a0022ffd14a003a3ea),
    .INIT_67(256'h022ffd14b00206a0022ffd14a00363ea022ffd14b0018bc0022ffd14a000bc02),
    .INIT_68(256'h022ffd14a00363d8022ffd0ba270d040022ffd14b0009002022ffd14a00206a0),
    .INIT_69(256'h022ffd14a001da20022ffd14b00323d8022ffd14a001fb00022ffd14b001da00),
    .INIT_6A(256'h022ffd2fb161fb00022ffd06b201da80022ffd0b216323d8022ffd14b001fb00),
    .INIT_6B(256'h022ffd20a25323d8022ffd0b92b1fb00022ffd0b82a1daa0022ffd00160323d8),
    .INIT_6C(256'h022ffd0ba251dae0022ffd01b00323d8022ffd20a4f1fb00022ffd20a311dac0),
    .INIT_6D(256'h022ffd14a001fb01022ffd0ba261da20022ffd14b00323d8022ffd14a0e1fb00),
    .INIT_6E(256'h022ffd14a00323d8022ffd14b001fb01022ffd14a001da80022ffd14b00323d8),
    .INIT_6F(256'h022ffd2f2191dac0022ffd062b0323d8022ffd0b2191fb01022ffd14b001daa0),
    .INIT_70(256'h022ffd14b001fb02022ffd14a001da00022ffd14b00323d8022ffd14a001fb01),
    .INIT_71(256'h022ffd14b00323d8022ffd14a001fb02022ffd14b001da20022ffd14a00323d8),
    .INIT_72(256'h022ffd14a001daa0022ffd0ba27323d8022ffd14b001fb02022ffd14a001da80),
    .INIT_73(256'h022ffd14a001fb02022ffd14b001dac0022ffd14a00323d8022ffd14b001fb02),
    .INIT_74(256'h022ffd2fb18323d8022ffd06b201fb03022ffd0b2181da00022ffd14b00323d8),
    .INIT_75(256'h022ffd20a25223ea022ffd0b92d323d8022ffd0b82c1fb03022ffd001501dae0),
    .INIT_76(256'h022ffd0ba25001b0022ffd01b00000a0022ffd20a4f20894022ffd20a31206da),
    .INIT_77(256'h022ffd14a0000bc0022ffd0ba26208e2022ffd14b00208b5022ffd14a0e208d2),
    .INIT_78(256'h022ffd14a00206b4022ffd14b0000ce0022ffd14a00206b4022ffd14b0000cf0),
    .INIT_79(256'h022ffd2f21b206b4022ffd062b000cb0022ffd0b21b206b4022ffd14b0000cd0),
    .INIT_7A(256'h022ffd14b0020779022ffd14a00206da022ffd14b00223ea022ffd14a00208a3),
    .INIT_7B(256'h022ffd14b0020894022ffd14a00206da022ffd14b0020716022ffd14a0022008),
    .INIT_7C(256'h022ffd14a002b40f022ffd0ba272b20f022ffd14b00208a3022ffd14a0020135),
    .INIT_7D(256'h022ffd14a0020779022ffd14b002074b022ffd14a0001002022ffd14b002b80f),
    .INIT_7E(256'h022ffd2fb1a20135022ffd06b2020894022ffd0b21a206da022ffd14b0022008),
    .INIT_7F(256'h022ffd20a252b80f02bff30b92f2b40f02bff00b82e2b20f022ffd00140208a3),
    .INITP_00(256'hd6f4e648c070fa75da61f9cad0d2f6d1f3f8fee45e6cec695a5b76e156f463c4),
    .INITP_01(256'hdc66e66f5bf4c67ac5eb7fe04de2e277dd6a5873cc76557dd263cd59dc61eae0),
    .INITP_02(256'h7cf5e76c747f7fe2d6e1ff4ce9fc41e57ecb71ec41e27eceeaea417b6d496a75),
    .INITP_03(256'h416cddc47963e9f1767078eff34efd74f9eb61f7fbff4fe5e5797f63746a61c8),
    .INITP_04(256'h706e6b66dbed74e4ec454fd273fed479d64e606bcae75cf2706dd177d1646270),
    .INITP_05(256'he27ce454f5e1f8fcc1d179eb684e4556547e42c7f160e5e0fc6179647b697576),
    .INITP_06(256'h60ffd1c85cf46b575d5eee4a6ad0766fe0c761cbf4e265f6ec6f6e6268707ef3),
    .INITP_07(256'h44c1645b64d9f655edcbf049db77d8dee773fcd863dae66b5d66f845c344fa47),
    .INITP_08(256'hf673d0dfc9c5554b5dc04f405fd159d8e9f5eff6c46ec9f05e6b45f6616341df),
    .INITP_09(256'hf54eda584d59cdc0d5c75aeacafedb69d5e35c56c7cd76cd66f647eeec47cc40),
    .INITP_0A(256'hc173d2417349e941f64170c94ceee9c8cfe1e1d156e5fac9dcfd597848794878),
    .INITP_0B(256'he8c0edfff963fd5ff0c2f5e2fd4655cedec1c1634e7b5b42d4e04bc5c9e5ccfb),
    .INITP_0C(256'hea53ecd6eac9ead24dc6c270567e426f506171c56ec34cf3f47e4bc56be6e649),
    .INITP_0D(256'h5947466641fdcf62def66247f04752f1f67e5fdcc5f0d97ec9625d60d5e4f8c9),
    .INITP_0E(256'hcc68764ee5d9537666e5c652c364c162d8e741fb4564fbcf62d8ea41fb4362de),
    .INITP_0F(256'h7b5b7c5d5c635a794eebceefd276fc457f436b5a6d43f2dfc04ec5eac6e9c660),
